* SPICE3 file created from inverter.ext - technology: scmos

.option scale=1u

M1000 out in vdd vdd pfet w=10 l=3
+  ad=110 pd=42 as=70 ps=34
M1001 out in gnd_ Gnd nfet w=8 l=3
+  ad=80 pd=36 as=56 ps=30
C0 vdd in 2.10fF
C1 gnd_ Gnd 4.89fF
C2 out Gnd 3.57fF
C3 in Gnd 8.54fF
